library ieee;
use ieee.std_logic_1164.all;
use std.env.stop;
use ieee.numeric_std.all;

library work;
use work.logger.all;
use work.ss_math.all;
use work.operations.all;

entity execute_tb is
end execute_tb;

architecture test of execute_tb is
	
	signal AluSrc			:	std_logic := '0';
	signal AluControl		:	std_logic_vector(3 downto 0) := (others => '0');
	signal PC_E, signImm_E		:	data_bus := (others => '0');
	signal readData1_E		:	data_bus := (others => '0');
	signal readData2_E		:	data_bus := (others => '0');
	signal PCBranch_E, aluResult_E	:	data_bus := (others => '0');
	signal writeData_E		:	data_bus := (others => '0');
	signal zero_E			:	std_logic := '0'
	
	constant DEC_500	:	data_bus := int_to_vec(500, data_bus'length);
	constant DEC_400	:	data_bus := int_to_vec(400, data_bus'length);
	constant DEC_200	:	data_bus := int_to_vec(200, data_bus'length);
	constant DEC_100	:	data_bus := int_to_vec(100, data_bus'length);

	type test_vector is record
		AluSrc			:	std_logic;
		AluControl		:	std_logic_vector(3 downto 0);
		PC_E, signImm_E		:	data_bus;
		readData1_E		:	data_bus;
		readData2_E		:	data_bus;
		PCBranch_E, aluResult_E	:	data_bus;
		writeData_E		:	data_bus;
		zero_E			:	std_logic;
	end record test_vector;

	type test_data is array (natural range <>) of test_vector;

	constant tests: test_data := (
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('1', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),
	('0', ADD_HEX, DEC_100, DEC_100, DEC_100, DEC_200, DEC_500, DEC_200, DEC_300, '0'),

	
begin
	dut : entity work.execute
	port map(AluSrc => AluSrc, AluControl => AluControl,
		PC_E => PC_E, signImm_E => signImm_E,
		readData1_E => readData1_E, readData2_E => readData2_E,
		PCBranch_E => PCBranch_E, aluResult_E => aluResult_E,
		writeData_E => writeData_E, zero_E => zero_E);

	stimulus : process
	begin
		wait for 10 ns;
		for i in tests'range loop
			AluSrc	<=	tests(i).AluSrc;
			AluControl	<= tests(i).AluControl;
			PC_E		<= tests(i).PC_E;
			signImm_E	<= tests(i).signImm_E;
			readData1_E	<= tests(i).readData1_E;
			readData2_E	<= tests(i).readData2_E;
			wait for 1 ns;
			checkEqual(PCBranh_E, tests(i).PCBranch_E, "Testing PC Branch");
			checkEqual(aluResult_E, tests(i).aluResult_E, "Testing PC Branch");
			checkEqual(writeData_E, tests(i).writeData_E, "Testing PC Branch");
			checkEqual(zero_E, tests(i).zero_E, "Testing PC Branch");
		end loop;		
			
	end process;
end architecture;
			
					
	
